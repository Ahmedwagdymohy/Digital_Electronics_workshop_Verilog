module full_adder_dataflow (A, B , CIN , CARRY, OUT );
// IN GALLERY
