module and_gateee (A,B,OUT);
input A,B;
output OUT;
assign OUT=A&B;
endmodule