module sync_reset(A,B,sel, clk, Q);
input A,B,clk,sel;
output reg Q;
always@(posedge CLK) begin
    if(sel)
    


end